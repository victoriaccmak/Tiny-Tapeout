/*
 * Copyright (c) 2024 Uri Shaked
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_vga_example(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,   // Dedicated outputs
  input  wire [7:0] uio_in,   // IOs: Input path
  output wire [7:0] uio_out,  // IOs: Output path
  output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
  input  wire       ena,      // always 1 when powered
  input  wire       clk,      // clock
  input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  wire [1:0] R;
  wire [1:0] G;
  wire [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;
  wire sound;

  // TinyVGA PMOD
  assign uo_out = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  assign uio_out = 0;
  assign uio_oe  = 0;
  wire _unused_ok = &{ena, ui_in, uio_in};

  reg [9:0] counter;

  hvsync_generator hvsync_gen(
    .clk(clk),
    .reset(~rst_n),
    .hsync(hsync),
    .vsync(vsync),
    .display_on(video_active),
    .hpos(pix_x),
    .vpos(pix_y)
  );

  // --- Dithering logic for color #522a1d ---
  wire dither = pix_x[0] ^ pix_y[0]; // simple 2x2 pattern

  wire [1:0] red_level   = dither ? 2'b10 : 2'b01; // alternate between 1 and 2
  wire [1:0] green_level = dither ? 2'b01 : 2'b00; // alternate between 0 and 1
  wire [1:0] blue_level  = 2'b00;                  // very low blue component

  assign R = video_active ? red_level   : 2'b00;
  assign G = video_active ? green_level : 2'b00;
  assign B = video_active ? blue_level  : 2'b00;

  always @(posedge vsync or negedge rst_n) begin
    if (~rst_n)
      counter <= 0;
    else
      counter <= counter + 1;
  end

endmodule
